LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY controle IS 
	PORT (
		F : IN STD_LOGIC_VECTOR(0 TO 2);
		EnA, EnB, InvA, InvB, C0, O1, O0 : OUT STD_LOGIC
	);
END controle;

ARCHITECTURE funccontrole OF controle IS

BEGIN
	
END funccontrole;